//                              -*- Mode: Verilog -*-
// Filename        : testbench.v
// Description     : VScale RiscV WV SoC Testbench
// Author          : Philip Tracton
// Created On      : Tue Dec  6 21:11:19 2016
// Last Modified By: Philip Tracton
// Last Modified On: Tue Dec  6 21:11:19 2016
// Update Count    : 0
// Status          : Unknown, Use with caution!


module testbench (/*AUTOARG*/ ) ;
   
endmodule // testbench
